//`include "LS_controller.sv"
//`include "Pipeline_reg.sv"
module Controller (
    input clk,
    input rst,
    stall,
    input logic [31:0] instruction,
    input logic br_taken,
    flush,
    gemm_done,
    output logic [3:0] ALUctrl,
    output logic mem_wr_ppl,
    mem_read_ppl,
    output logic A_sel,
    B_sel,
    reg_wr_ppl,
    PC_sel_ppl,
    is_mret_ppl,
    csr_reg_r_ppl,
    csr_reg_wr_ppl,
    //gemm signals
    is_GemmInstr_ppl,
    output logic [1:0] wb_sel_ppl
);
  localparam R_type = 5'b01100;
  localparam I_type = 5'b00100;
  localparam Load_type = 5'b00000;
  localparam S_type = 5'b01000;
  localparam B_type = 5'b11000;
  localparam JAL_TYPE = 5'b11011;
  localparam Jalr_type = 5'b11001;
  localparam lui_type = 5'b01101;
  localparam auipc_type = 5'b00101;
  localparam csr_type = 5'b11100;
  localparam GEMM_type = 5'b000010;
  logic [6:0] opcode;
  logic func7, func7_mret, is_mret, csr_reg_r, csr_reg_wr;
  logic [2:0] func3;
  assign func3 = instruction[14:12];
  assign opcode = instruction[6:0];
  assign func7 = instruction[30];
  assign func7_mret = instruction[29];
  logic [1:0] wb_sel;
  logic PC_sel, reg_wr, mem_wr, mem_read;
  logic is_GemmInstr;
  // mul     rd rs1 rs2 31..25=1 14..12=0 6..2=0x0C 1..0=3
  // add     rd rs1 rs2 31..25=0  14..12=0 6..2=0x0C 1..0=3
  // sub     rd rs1 rs2 31..25=32 14..12=0 6..2=0x0C 1..0=3
  // sll     rd rs1 rs2 31..25=0  14..12=1 6..2=0x0C 1..0=3
  // slt     rd rs1 rs2 31..25=0  14..12=2 6..2=0x0C 1..0=3
  // sltu    rd rs1 rs2 31..25=0  14..12=3 6..2=0x0C 1..0=3
  // xor     rd rs1 rs2 31..25=0  14..12=4 6..2=0x0C 1..0=3
  // srl     rd rs1 rs2 31..25=0  14..12=5 6..2=0x0C 1..0=3
  // sra     rd rs1 rs2 31..25=32 14..12=5 6..2=0x0C 1..0=3
  // or      rd rs1 rs2 31..25=0  14..12=6 6..2=0x0C 1..0=3
  // and     rd rs1 rs2 31..25=0  14..12=7 6..2=0x0C 1..0=3
  always_comb begin
    case (opcode[6:2])
      R_type: begin
        casez ({
          instruction[25], instruction[30], func3
        })
          5'b00000: ALUctrl = 4'd0;  //ADD
          5'b01000: ALUctrl = 4'd1;  //Sub
          5'b00001: ALUctrl = 4'd2;  //SLL
          5'b00010: ALUctrl = 4'd3;  //SLT
          5'b00100: ALUctrl = 4'd4;  //XOR
          5'b00011: ALUctrl = 4'd5;  //SLTU
          5'b00101: ALUctrl = 4'd6;  //SRL
          5'b01101: ALUctrl = 4'd7;  //SRA
          5'b00110: ALUctrl = 4'd8;  //OR
          5'b00111: ALUctrl = 4'd9;  //AND
          5'b10000: ALUctrl = 4'd11;  //MUL
          5'b10001: ALUctrl = 4'd12;  //MULH
          5'b10010: ALUctrl = 4'd13;  //MULHSU
          5'b10011: ALUctrl = 4'd14;  //MULHU
          default:  ALUctrl = 4'bXXXX;
        endcase
        A_sel = 1;
        PC_sel = 0;
        mem_wr = 0;
        mem_read = '0;
        B_sel = 0;
        wb_sel = 2'b01;
        reg_wr = 1;
        csr_reg_r = 1'b0;
        csr_reg_wr = 1'b0;
        is_mret = 1'b0;
        is_GemmInstr = 1'b0;
      end
      I_type: begin
        casez ({
          func7, func3
        })
          4'b?000: ALUctrl = 4'd0;  //ADD
          4'b?001: ALUctrl = 4'd2;  //SLL
          4'b?010: ALUctrl = 4'd3;  //SLT
          4'b?100: ALUctrl = 4'd4;  //XOR
          4'b?011: ALUctrl = 4'd5;  //SLTU
          4'b0101: ALUctrl = 4'd6;  //SRL
          4'b1101: ALUctrl = 4'd7;  //SRA
          4'b?110: ALUctrl = 4'd8;  //OR
          4'b?111: ALUctrl = 4'd9;  //AND
          default: begin
            ALUctrl = 4'bXXXX;
          end
        endcase
        mem_wr = 0;
        mem_read = '0;
        A_sel = 1;
        PC_sel = 0;
        B_sel = 1;
        wb_sel = 2'b01;
        reg_wr = 1;
        csr_reg_r = 1'b0;
        csr_reg_wr = 1'b0;
        is_mret = 1'b0;
        is_GemmInstr = 1'b0;
      end
      Load_type: begin
        mem_wr = 0;
        mem_read = 1'b1;
        A_sel = 1;
        PC_sel = 0;
        B_sel = 1;
        wb_sel = 2'b10;
        reg_wr = 1;
        ALUctrl = 4'd0;
        csr_reg_r = 1'b0;
        csr_reg_wr = 1'b0;
        is_mret = 1'b0;
        is_GemmInstr = 1'b0;
      end
      S_type: begin
        mem_wr = 1;
        mem_read = '0;
        A_sel = 1;
        PC_sel = 0;
        B_sel = 1;
        wb_sel = 'x;
        reg_wr = 0;
        ALUctrl = 4'd0;
        csr_reg_r = 1'b0;
        csr_reg_wr = 1'b0;
        is_mret = 1'b0;
        is_GemmInstr = 1'b0;
      end
      B_type: begin
        mem_wr = 0;
        mem_read = '0;
        A_sel = 0;
        B_sel = 1;
        wb_sel = 'x;
        reg_wr = 0;
        ALUctrl = 4'd0;
        csr_reg_r = 1'b0;
        csr_reg_wr = 1'b0;
        is_mret = 1'b0;
        is_GemmInstr = 1'b0;
        case (br_taken)
          0: PC_sel = 0;
          1: PC_sel = 1;
          default: PC_sel = 'x;
        endcase
      end
      JAL_TYPE: begin
        mem_wr = 0;
        mem_read = '0;
        A_sel = 0;
        B_sel = 1;
        // wb_sel = 2'b00;
        wb_sel = 2'b00;
        // reg_wr = 1;
        reg_wr = 1'b1;
        ALUctrl = 4'd0;
        PC_sel = 1'b1;
        csr_reg_r = 1'b0;
        csr_reg_wr = 1'b0;
        is_mret = 1'b0;
        is_GemmInstr = 1'b0;
      end
      Jalr_type: begin
        mem_wr = 0;
        mem_read = '0;
        A_sel = 1;
        B_sel = 1;
        wb_sel = 2'b00;
        reg_wr = 1'b1;
        ALUctrl = 4'd0;
        PC_sel = 1'b1;
        csr_reg_r = 1'b0;
        csr_reg_wr = 1'b0;
        is_mret = 1'b0;
        is_GemmInstr = 1'b0;
      end
      lui_type: begin
        mem_wr = 0;
        mem_read = '0;
        A_sel = 1'bx;
        B_sel = 1;
        wb_sel = 2'b01;
        reg_wr = 1'b1;
        ALUctrl = 4'd10;
        PC_sel = 1'b0;
        csr_reg_r = 1'b0;
        csr_reg_wr = 1'b0;
        is_mret = 1'b0;
        is_GemmInstr = 1'b0;
      end
      auipc_type: begin
        mem_wr = 0;
        mem_read = '0;
        A_sel = 0;
        B_sel = 1;
        wb_sel = 2'b01;
        reg_wr = 1;
        ALUctrl = 4'd0;
        PC_sel = 1'b0;
        csr_reg_r = 1'b0;
        csr_reg_wr = 1'b0;
        is_mret = 1'b0;
        is_GemmInstr = 1'b0;
      end
      csr_type: begin
        mem_wr = 0;
        mem_read = '0;
        A_sel = 1;
        B_sel = 1'bx;
        wb_sel = 2'b11;
        reg_wr = 1'b1;
        ALUctrl = 4'd0;
        PC_sel = 1'b0;
        is_GemmInstr = 1'b0;
        casez ({
          func7_mret, func3
        })
          4'b1000: begin
            csr_reg_r = 1'b0;
            csr_reg_wr = 1'b0;
            is_mret = 1'b1;
          end
          4'b?001: begin
            csr_reg_r = 1'b1;
            csr_reg_wr = 1'b1;
            is_mret = 1'b0;
          end
          default: begin
            csr_reg_r = 1'b0;
            csr_reg_wr = 1'b0;
            is_mret = 1'b0;
          end
        endcase
      end
      GEMM_type: begin
        ALUctrl = 4'bXXXX;
        A_sel = 1;
        B_sel = 0;
        PC_sel = 0;
        mem_wr = 0;
        mem_read = '0;
        wb_sel = 2'b01;
        reg_wr = 1'b0;
        csr_reg_r = 1'b0;
        csr_reg_wr = 1'b0;
        is_mret = 1'b0;
        is_GemmInstr = 1'b1;
      end
      default: begin
        mem_wr = 'x;
        mem_read = 'x;
        B_sel = 'x;
        A_sel = 'x;
        wb_sel = 'x;
        reg_wr = 'x;
        ALUctrl = 'x;
        PC_sel = 'x;
        csr_reg_r = 1'bx;
        csr_reg_wr = 1'bx;
        is_mret = 1'bx;
        is_GemmInstr = 1'b0;
      end
    endcase
  end
  // 
  Pipeline_reg #(
      .WIDTH(1),
      .reset(0)
  ) Pipeline1 (
      .clk(clk),
      .flush(flush),
      .stall(stall),
      .in(reg_wr),
      .out(reg_wr_ppl)
  );
  Pipeline_reg #(
      .WIDTH(1),
      .reset(0)
  ) pipeline2 (
      .clk(clk),
      .flush(flush),
      .stall(stall),
      .in(mem_wr),
      .out(mem_wr_ppl)
  );
  Pipeline_reg #(
      .WIDTH(2),
      .reset(0)
  ) pipeline3 (
      .clk(clk),
      .flush(flush),
      .stall(stall),
      .in(wb_sel),
      .out(wb_sel_ppl)
  );

  Pipeline_reg #(
      .WIDTH(1),
      .reset(0)
  ) Pipieline4 (
      .clk(clk),
      .flush(flush),
      .stall(stall),
      .in(PC_sel),
      .out(PC_sel_ppl)
  );
  Pipeline_reg #(
      .WIDTH(1),
      .reset(0)
  ) Pipeline_reg_instance (
      .clk(clk),
      .flush(flush),
      .stall(stall),
      .in(mem_read),
      .out(mem_read_ppl)
  );
  Pipeline_reg #(
      .WIDTH(1),
      .reset(0)
  ) Pipeline_ismret (
      .clk(clk),
      .flush(flush),
      .stall(stall),
      .in(is_mret),
      .out(is_mret_ppl)
  );
  Pipeline_reg #(
      .WIDTH(1),
      .reset(0)
  ) Pipeline_csr_reg_r (
      .clk(clk),
      .flush(flush),
      .stall(stall),
      .in(csr_reg_r),
      .out(csr_reg_r_ppl)
  );
  Pipeline_reg #(
      .WIDTH(1),
      .reset(0)
  ) Pipeline_csr_reg_wr (
      .clk(clk),
      .flush(flush),
      .stall(stall),
      .in(csr_reg_wr),
      .out(csr_reg_wr_ppl)
  );

  Pipeline_reg #(
      .WIDTH(1),
      .reset(0)
  ) Pipeline_reg_instance1 (
      .clk(clk),
      .flush(flush),
      .stall(stall),
      .in(is_GemmInstr),
      .out(is_GemmInstr_ppl)
  );
endmodule
